`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   15:03:13 02/07/2018
// Design Name:   rippler
// Module Name:   /media/raditya/822A-B6CA/CS220Labs/Lab3_2/ripple_led/rippler_top.v
// Project Name:  ripple_led
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: rippler
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module rippler_top;

	// Inputs
	reg clk;

	// Outputs
	wire led0;
	wire led1;
	wire led2;
	wire led3;
	wire led4;
	wire led5;
	wire led6;
	wire led7;

	// Instantiate the Unit Under Test (UUT)
	rippler uut (
		.clk(clk), 
		.led0(led0), 
		.led1(led1), 
		.led2(led2), 
		.led3(led3), 
		.led4(led4), 
		.led5(led5), 
		.led6(led6), 
		.led7(led7)
	);

	always @(led0) begin
		$display("time=%d: clk=%b, led0=%b, led1=%b, led2=%b, led3=%b, led4=%b, led5=%b, led6=%b, led7=%b", $time, clk, led0, led1, led2, led3, led4, led5, led6, led7);
   end

   initial begin
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		clk=0;
      #5
      clk=1;
      #5
		$finish;
	end

endmodule

